package wifii_pkg;

endpackage
